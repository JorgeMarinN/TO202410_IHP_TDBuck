** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/tb_LSHL_v3p1.sch
**.subckt tb_LSHL_v3p1
VCC VCC GND 1.2
VSS VSS GND 0
VIN VIN VSS PULSE(0 3.3 3u 100p 100p 12u 24u)
C1 VOUT VSS 10f m=1
X1 VIN VOUT VCC VSS LSHL_v3p1
VCC1 VH GND 3.3
**** begin user architecture code


.option scale=1e-6
.save v(vin) v(vout)
.control
tran 100p 6u
plot v(vin) v(vout)
plot v(vin) v(vout)+2
.endc

.measure tran tdelay
+ TRIG tran1.V(VIN) TD=0u VAL=0.6 RISE=1
+ TARG tran1.V(VOUT) TD=0u VAL=0.6 RISE=1






.param corner=0

.if (corner==0)
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.endif

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  /home/designer/shared/TO202410_IHP_TDBuck/xschem/LSHL_v3p1.sym # of pins=4
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/LSHL_v3p1.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/LSHL_v3p1.sch
.subckt LSHL_v3p1 Vs Vg VDIG VSS
*.iopin VDIG
*.ipin Vs
*.opin Vg
*.iopin VSS
XMD5 VgMD2 Vs VDIG VDIG sg13_hv_pmos w=1u l=0.4u ng=1 m=2
XMD6 VgMD2 Vs VSS VSS sg13_hv_nmos w=1u l=0.45u ng=1 m=1
x7 net1 VDIG VSS Vg sg13g2_buf_4
x1 VgMD2 VDIG VSS net1 sg13g2_inv_1
.ends

.GLOBAL GND
.end
