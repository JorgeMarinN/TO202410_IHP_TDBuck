** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/inv_VCO_nmoshv.sch
.subckt inv_VCO_nmoshv D S G B
*.PININFO D:B S:B G:B B:B
M1 D G net1 B sg13_hv_nmos l=5u w=2u ng=1 m=1
.ends
.end
