** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/TB_DCDCBuck_GateDrivers_NOL.sch
**.subckt TB_DCDCBuck_GateDrivers_NOL
X1 Vg_M1 Vg_M2 net1 net6 Vo DCDC_Buck
Vdd Vdd GND {Vdd}
Vg1 Vs GND PULSE(0 {Vdd} 0 {TR} {TF} {T*D} {T} 0)
V_Iin VH net1 0
.save i(v_iin)
X2 Vs_M1 Vg_M1 net2 net3 GND GateDriver
X3 Vs_M2 Vg_M2 net4 net5 GND GateDriver
Vdd1 VH GND {VH}
V_Igd_VH1 VH2 net3 0
.save i(v_igd_vh1)
V_Igd_VH2 VH2 net5 0
.save i(v_igd_vh2)
V_Igd_Vdd2 Vdd net4 0
.save i(v_igd_vdd2)
V_Igd_Vdd1 Vdd net2 0
.save i(v_igd_vdd1)
Vdd2 Vdd2 GND {Vdd}
Vdd3 VH2 GND {VH}
x4 Vdd2 GND Vs_M1 Vs Vs_M2 NOL_v2p2_AM
**** begin user architecture code


*M1 hvPMOS
.param temp=27
.param mult_M1 = 12000
.param w_M1 =10u
.param l_M1 = 0.4u
.param ng_M1 = 1

*M2 hvNMOS
.param mult_M2 = 4000
.param w_M2 =10u
.param l_M2 =0.45u
.param ng_M2 =1








.param Vdd = 1.2
.param VH = 3.3
.param Del = 0

*.param D = 0.42
*.param T = 1u
*.param TR = 7n
*.param TF = 7n
*.param TdR = 0.1u
*.param TdF = 0.1u

*.param D = 0.6364
.param D = 0.615
.param T = 0.1u
.param TR = 1n
.param TF = 1n
.param TdR = 1.5n
.param TdF = 1.5n
*.param TdR = 1n
*.param TdF = 1n


.param temp = 27





*Parametros
*Filtro
*.param L = 1.37u
*.param R = 0.9
*.param C = 416n

* Io=2A 10MHz
*.param L = 137.5n
*.param R = 0.6
*.param C = 62.5n

* Io=1A 10MHz
*.param L = 275n
*.param R = 1.2
*.param C = 31.25n

* Io=1A 10MHz
.param L = 1u
.param R = 1.2
.param C = 1u





*.save all
.save v(vo)
+ @n.x1.xm1.nsg13_hv_pmos[ids]
+ @n.x1.xm2.nsg13_hv_nmos[ids]
.param SimTime = 5u

.option method=gear

.control
reset
set color0 = white
tran 100p 5u
let Io = i(v.x1.V_Io)
let Id_M1 = @n.x1.xm1.nsg13_hv_pmos[ids]
let Id_M2 = @n.x1.xm2.nsg13_hv_nmos[ids]
let Po = Io*v(Vo)
let I_in = i(V_Iin)
let Pin = I_in*v(VH)
let Vsd_M1 = v(VH) - v(x1.Vc)
let Vds_M2 = v(x1.Vc)
let P_M1 = Vsd_M1*Id_M1
let P_M2 = -Vds_M2*Id_M2
let P_GD_Vdd = v(Vdd)*(i(V_Igd_Vdd1)+i(V_Igd_Vdd2))
let P_GD_VH = v(VH)*(i(V_Igd_VH1)+i(V_Igd_VH2))
let DataMeasBegin = SimTime-1u

meas tran Vo_mean AVG v(Vo) from=4u to=5u
meas tran Io_mean AVG Io from=4u to=5u
meas tran Po_mean AVG Po from=4u to=5u
meas tran Pin_mean AVG Pin from=4u to=5u
meas tran P_M1_mean AVG P_M1 from=4u to=5u
meas tran P_M2_mean AVG P_M2 from=4u to=5u
meas tran P_GD_Vdd_mean AVG P_GD_Vdd from=4u to=5u
meas tran P_GD_VH_mean AVG P_GD_VH from=4u to=5u

let P_GD = P_GD_Vdd_mean+P_GD_VH_mean
let Pin_tot_mean = P_GD + Pin_mean
let eff = 100*Po_mean/Pin_tot_mean
let eff_DCDC = 100*Po_mean/Pin_mean
let loss_M1 = 100*P_M1_mean/Pin_tot_mean
let loss_M2 = 100*P_M2_mean/Pin_tot_mean
let loss_GD = 100*P_GD/Pin_tot_mean
let sumaPot = eff+loss_M1+loss_M2+loss_GD
print eff eff_DCDC loss_M1 loss_M2 loss_GD sumaPot

plot Io i(v.x1.V_IL)
plot Id_M1 Id_M2
plot v(Vo)
plot Po Pin
*plot P_M1 P_M2
plot v(x1.Vc)
plot v(Vg_M1) v(Vg_M2)
.endc



.end




.param temp=27

*.param mult_13 = 1
*.param mult_24 = 6
*.param mult_5 = 100
*.param mult_6 = 100
*.param mult_7 = 200
*.param mult_8 = 200
*.param mult_9 = 5
*.param mult_10 = 5

.param mult_13 = 1
.param mult_24 = 6
*.param mult_5 = 25
*.param mult_6 = 25
.param mult_5 = 30
.param mult_6 = 25
.param mult_7 = 250
.param mult_8 = 200
*.param mult_7 = 75
*.param mult_8 = 60
.param mult_9 = 15
.param mult_10 = 15

.param ng_13 = 1
.param ng_24 = 1
.param ng_5 = 1
.param ng_6 = 1
.param ng_7 = 1
.param ng_8 = 1
.param ng_9 = 1
.param ng_10 = 1

.param l_1357 = 0.4u
*.param w_1357 = 0.3u
.param w_1357 = 10u
.param l_2468 = 0.45u
*.param w_2468 = 0.3u
.param w_2468 = 10u
.param l_9 = 0.13u
.param w_9 = 0.15u
.param l_10 = 0.13u
.param w_10 = 0.15u





.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.lib cornerMOShv.lib mos_tt
.lib cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ




**** end user architecture code
**.ends

* expanding   symbol:  DCDC_Buck.sym # of pins=5
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/DCDC_Buck.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/DCDC_Buck.sch
.subckt DCDC_Buck VgM1 VgM2 Vin GND Vo
*.iopin Vin
*.ipin VgM1
*.ipin VgM2
*.iopin Vo
*.iopin GND
XM2 Vc VgM2 GND GND sg13_hv_nmos w={w_M2} l={l_M2} ng={ng_M2} m={mult_M2}
XM1 Vc VgM1 Vin Vin sg13_hv_pmos w={w_M1} l={l_M1} ng={ng_M1} m={mult_M1}
L1 net2 net1 {L} m=1
C1 net1 GND {C} m=1
V_Io net1 Vo 0
.save i(v_io)
V_IL Vc net2 0
.save i(v_il)
R1 Vo GND {R} m=1
.ends


* expanding   symbol:  GateDriver.sym # of pins=5
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/GateDriver.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/GateDriver.sch
.subckt GateDriver Vs Vg Vdd VH GND
*.iopin VH
*.iopin Vdd
*.ipin Vs
*.opin Vg
*.iopin GND
XMD9 VgMD2 Vs Vdd Vdd sg13_lv_pmos w={w_9} l={l_9} ng={ng_9} m={mult_9}
XMD10 VgMD2 Vs GND GND sg13_lv_nmos w={w_10} l={l_10} ng={ng_10} m={mult_10}
XMD1 VgMD5 net1 VH VH sg13_hv_pmos w={w_1357} l={l_1357} ng={ng_13} m={mult_13}
XMD3 net1 VgMD5 VH VH sg13_hv_pmos w={w_1357} l={l_1357} ng={ng_13} m={mult_13}
XMD5 net2 VgMD5 VH VH sg13_hv_pmos w={w_1357} l={l_1357} ng={ng_5} m={mult_5}
XMD7 Vg VgMd78 VH VH sg13_hv_pmos w={w_1357} l={l_1357} ng={ng_7} m={mult_7}
XMD2 VgMD5 VgMD2 GND GND sg13_hv_nmos w={w_2468} l={l_2468} ng={ng_24} m={mult_24}
XMD4 net1 Vs GND GND sg13_hv_nmos w={w_2468} l={l_2468} ng={ng_24} m={mult_24}
XMD6 net2 Vs GND GND sg13_hv_nmos w={w_2468} l={l_2468} ng={ng_6} m={mult_6}
XMD8 Vg VgMd78 GND GND sg13_hv_nmos w={w_2468} l={l_2468} ng={ng_8} m={mult_8}
VIg78 net2 VgMd78 0
.save i(vig78)
.ends


* expanding   symbol:  NOL_v2p2_AM.sym # of pins=5
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/NOL_v2p2_AM.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/NOL_v2p2_AM.sch
.subckt NOL_v2p2_AM VCC VSS VCP CLK VCN
*.iopin CLK
*.iopin VCP
*.iopin VCN
*.iopin VCC
*.iopin VSS
x5 CLK VCC VSS A1 sg13g2_inv_1
x3 A1 B1 VCC VSS C1 sg13g2_nor2_1
x1 B2 CLK VCC VSS C2 sg13g2_nor2_1
x2 B1 VCC VSS net1 sg13g2_inv_1
x6 B2 VCC VSS net2 sg13g2_inv_2
x7 net1 VCC VSS net3 sg13g2_inv_2
x8 net2 VCC VSS VCN sg13g2_inv_4
x9 net3 VCC VSS VCP sg13g2_inv_4
x11 VCC VSS C1 B2 delayRC2ns_v1p1
x4 VCC VSS C2 B1 delayRC2ns_v1p1
.ends


* expanding   symbol:  delayRC2ns_v1p1.sym # of pins=4
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/delayRC2ns_v1p1.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/delayRC2ns_v1p1.sch
.subckt delayRC2ns_v1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1 VIN VCC VSS net1 sg13g2_dlygate4sd3_1
x2 net1 VCC VSS VOUT sg13g2_dlygate4sd3_1
C1 net1 VSS 0.15p m=1
C2 VOUT VSS 0.15p m=1
.ends

.GLOBAL GND
.end
