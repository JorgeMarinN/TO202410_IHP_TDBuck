** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/tb_NOL_vto1p1.sch
**.subckt tb_NOL_vto1p1
VCC VCC GND 1.2
VSS VSS GND 0
VIN VIN VSS PULSE(0 1.2 25n 1p 1p 100n 200n)
C1 VCP VSS 10f m=1
C2 VCN VSS 10f m=1
x1 VCC VSS VCP VIN VCN NOL_vto1p1
**** begin user architecture code


.save v(vin) v(vcp) v(vcn)
.control
tran 100p 300n
plot v(vin) v(vcp) v(vcn)
plot v(vin) v(vcp)+1.5 v(vcn)+3
.endc

.measure tran tdead_fall
+ TRIG tran1.V(vcn) TD=0u VAL=0.6 FALL=1
+ TARG tran1.V(vcp) TD=0u VAL=0.6 FALL=1


.measure tran tdead_rise
+ TRIG tran1.V(vcp) TD=0u VAL=0.6 RISE=1
+ TARG tran1.V(vcn) TD=0u VAL=0.6 RISE=1






.param corner=0

.if (corner==0)
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.endif

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  NOL_vto1p1.sym # of pins=5
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/NOL_vto1p1.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/NOL_vto1p1.sch
.subckt NOL_vto1p1 VCC VSS VCP CLK VCN
*.iopin CLK
*.iopin VCP
*.iopin VCN
*.iopin VCC
*.iopin VSS
x5 CLK VCC VSS A1 sg13g2_inv_1
x3 A1 B1 VCC VSS C1 sg13g2_nor2_1
x1 B2 CLK VCC VSS C2 sg13g2_nor2_1
x2 B1 VCC VSS net1 sg13g2_inv_1
x6 B2 VCC VSS net2 sg13g2_inv_2
x7 net1 VCC VSS net3 sg13g2_inv_2
x8 net2 VCC VSS VCN sg13g2_inv_4
x9 net3 VCC VSS VCP sg13g2_inv_4
x10 VCC VSS C1 B2 large_delay_vto1p1
x4 VCC VSS C2 B1 large_delay_vto1p1
.ends


* expanding   symbol:  large_delay_vto1p1.sym # of pins=4
** sym_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/large_delay_vto1p1.sym
** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1[0] VIN VCC VSS n2 sg13g2_dlygate4sd3_1
x1[1] n2 VCC VSS n3 sg13g2_dlygate4sd3_1
x1[2] n3 VCC VSS n4 sg13g2_dlygate4sd3_1
x1[3] n4 VCC VSS n5 sg13g2_dlygate4sd3_1
x1[4] n5 VCC VSS VOUT sg13g2_dlygate4sd3_1
.ends

.GLOBAL GND
.end
