** sch_path: /home/designer/shared/TO202410_IHP_TDBuck/xschem/VCDL_v3p1.sch
**.subckt VCDL_v3p1 VDD VCONT VOUT VIN VSS
*.ipin VIN
*.opin VOUT
*.iopin VDD
*.iopin VSS
*.ipin VCONT
XM9 net4 net4 VSS VSS sg13_hv_nmos w=5u l=0.5u ng=1 m=1
XM3 net3 net4 VSS VSS sg13_hv_nmos w=5u l=0.5u ng=1 m=1
XM5 net2 net4 VSS VSS sg13_hv_nmos w=3u l=0.5u ng=1 m=1
XM8 net4 VCONT VDD VDD sg13_hv_pmos w=4.5u l=7u ng=1 m=1
XM4 net3 net3 VDD VDD sg13_hv_pmos w=8u l=4u ng=1 m=1
XM6 net1 net3 VDD VDD sg13_hv_pmos w=5u l=4u ng=1 m=1
XM2 VOUT VIN net1 VDD sg13_hv_pmos w=2.5u l=5u ng=1 m=1
XM1 VOUT VIN net2 VSS sg13_hv_nmos w=1u l=5u ng=1 m=2
XM7 net4 VDD VDD VDD sg13_hv_pmos w=0.5u l=7u ng=1 m=1
**.ends
.end
