** sch_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/tb_PD_vto1p1.sch
**.subckt tb_PD_vto1p1
VCC Vdd GND {Vdd}
VSS Vss GND 0
Vg1 VIN_1 VSS PULSE(0 {Vdd} 0 {TR} {TF} {T*D} {T} 0)
C1 V_PWM Vss 1f m=1
Vg3 VIN_2 VSS PULSE(0 {Vdd} {Td} {TR} {TF} {T*D} {T} 0)
x1 Vdd Vss VIN_2 V_PWM VIN_1 PD_vto1p1
Vg2 Vctrl VSS PULSE(0 {Vdd} 0 {TR} {TF} {T*0.615} {T} 0)
**** begin user architecture code


.param corner=0

.if (corner==0)
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.endif

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param Vdd = 1.2
.param VH = 3.3
.param Del = 0

.param T = 0.1u
.param TR = 1p
.param TF = 1p
.param DD = 0.615

*Caso 1 - No funciona bien
*.param D = 0.8
*.param Td = 0.03u

*Caso 2 - Funciona bien
.param D = 0.5
.param Td = DD*T

*Caso 3 - Funciona bien
*.param D = 0.615
*.param Td = 0.03u

*Caso 4 - No funciona bien
*.param D = 0.615
*.param Td = 0.08u




.param temp = 27





.save all

.control
set color0 = white
tran 100p 300n
plot v(VIN_1) v(VIN_2)+1.5 v(V_PWM)+3
plot v(V_PWM) v(Vctrl)+1.5
.endc

*.measure tran tdead_fall
*+ TRIG tran1.V(vcn) TD=0u VAL=0.6 FALL=1
*+ TARG tran1.V(vcp) TD=0u VAL=0.6 FALL=1

*.measure tran t_large_delay
*+ TRIG tran1.V(x1.C1) TD=0u VAL=0.6 RISE=1
*+ TARG tran1.V(x1.B2) TD=0u VAL=0.6 RISE=1



**** end user architecture code
**.ends

* expanding   symbol:  PD_vto1p1.sym # of pins=5
** sym_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/PD_vto1p1.sym
** sch_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/PD_vto1p1.sch
.subckt PD_vto1p1 VCC VSS VINS V_PWM VINR
*.iopin V_PWM
*.iopin VCC
*.iopin VSS
*.iopin VINS
*.iopin VINR
x3 net2 V_PWM VCC VSS V_N sg13g2_nor2_1
x1 V_N net1 VCC VSS V_PWM sg13g2_nor2_1
x2 VCC VSS VFE1 VINR net2 SPG_vto1p1
x4 VCC VSS VFE1 VINS net1 SPG_vto1p1
.ends


* expanding   symbol:  ../SPG/SPG_vto1p1.sym # of pins=5
** sym_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/SPG/SPG_vto1p1.sym
** sch_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/SPG/SPG_vto1p1.sch
.subckt SPG_vto1p1 VCC VSS VFE VIN VRE
*.iopin VIN
*.iopin VFE
*.iopin VRE
*.iopin VCC
*.iopin VSS
x1 dly7 VCC VSS dly8 sg13g2_inv_1
x2 predly VCC VSS net2 sg13g2_inv_1
x3 net3 VCC VSS predly sg13g2_inv_1
x4 dly8 VCC VSS net1 sg13g2_inv_1
x5 VIN VCC VSS net3 sg13g2_inv_2
x6 predly VCC VSS V_gatein sg13g2_inv_8
x7 net2 dly8 VCC VSS VFE sg13g2_and2_2
x8 net1 predly VCC VSS VRE sg13g2_and2_2
x9 VCC VSS V_gatein dly7 large_delay_vto1p1
.ends


* expanding   symbol:  ../large_delay/large_delay_vto1p1.sym # of pins=4
** sym_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/large_delay/large_delay_vto1p1.sym
** sch_path: /home/designer/shared/TORepo_IHPNov2024_TDBuck/design_data/xschem/large_delay/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1[0] VIN VCC VSS n2 sg13g2_dlygate4sd3_1
x1[1] n2 VCC VSS n3 sg13g2_dlygate4sd3_1
x1[2] n3 VCC VSS n4 sg13g2_dlygate4sd3_1
x1[3] n4 VCC VSS n5 sg13g2_dlygate4sd3_1
x1[4] n5 VCC VSS VOUT sg13g2_dlygate4sd3_1
.ends

.GLOBAL GND
.end
